package packaga_alu;
  `include "transaction_alu.sv";
  `include "generator_alu.sv";
  `include "driver.sv";
  `include "monitor_alu.sv";
  `include "reference_model_alu.sv";
  `include "scoreboard_alu.sv";
  `include "environment_alu.sv";
  `include "test_alu.sv";
endpackage

