
package alu_pkg;
  `include "transaction_alu.sv"
  `include "generator_alu.sv"
  `include "driver_2.sv"
  `include "monitor_2.sv"
  `include "reference_model_alu.sv"
  `include "scoreboard_alu.sv"
  `include "environment_alu.sv"
  `include "test_alu.sv"
endpackage


