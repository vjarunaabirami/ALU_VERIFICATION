`define WIDTH 8
`define no_of_trans 30
